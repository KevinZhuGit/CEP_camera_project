`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 08/20/2022 09:57:31 PM
// Design Name: 
// Module Name: exp_ro_merge_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module exp_ro_merge_tb(

    );

	reg clk_100; initial clk_100 = 1'b0; always #5   clk_100 = ~clk_100; 
    reg clk_200; initial clk_200 = 1'b0; always #2.5 clk_200 = ~clk_200; 
    reg clk_7  ; initial clk_7   = 1'b0; always #35  clk_7   = ~clk_7; 
    wire CLKMi, TX_CLKi, TX_CLKi2;
    assign CLKMi = clk_100;
    assign TX_CLKi  = clk_100;
    assign TX_CLKi2 = clk_200;
    reg rst;

    wire [8:0] ROWADD;
    wire [8:0] ROWADD_EXP;
    wire [8:0] ROWADD_RO;
    
    wire ex_trigger;	
    wire re_busy;
    reg [31:0] wirerst, Select;


    // Readout
    parameter 
    	NUMROW_RO = 10,
    //T6 RO----------------------------------------
    	NUM_SAMP	= 2,
    	NUM_ROW		= 10,
    	T_PIX		= 100,
    	T1          = 5,
    	T2          = 100,
    	T3          = 20,
    	T4          = 10,
    	T5          = 14,
    	T6          = 6,
    	T7          = 17,
    	T8          = 14,
        TADC        = 13,
        TOSR        = 115,
        TReadRst    = 100,
        Tbuck       = 1652,
        T6_NUM_ADC_BITS = 14;
    // T7 RO----------------------------------------
     parameter  
        ADC1_Tcolumn           = 700,
    	ADC1_T1                = 10,
    	ADC1_T2_1              = 400,
    	ADC1_T2_0              = 420,
    	ADC1_T3                = 20*12,
    	ADC1_T4                = ADC1_T3+2,
    	ADC1_T5                = 4,
    	ADC1_T6                = 1,
    	ADC1_T7                = 22,
    	ADC1_T8                = 2,
    	ADC1_T9                = ADC1_T8+20,
    	ADC1_TADC              = 22,
    	ADC1_NUM_ROW           = NUMROW_RO,
    	ADC1_NUM_ADC_BITS      = 12,
    	ADC1_Wait              = 1024; 
    parameter
        ADC2_Tcolumn           = 36,
    	ADC2_T1                = 6,
    	ADC2_T2_1              = 0,
    	ADC2_T2_0              = 3,
    	ADC2_T3                = 0,
    	ADC2_T4                = 1,
    	ADC2_T5                = 1,
    	ADC2_T6                = 1,
    	ADC2_T7                = 11,
    	ADC2_T8                = 3,
    	ADC2_T9                = ADC2_T8+8,
    	ADC2_TADC              = 12,
    	ADC2_NUM_ROW           = NUMROW_RO,
    	ADC2_NUM_ADC_BITS      = 12,
    	ADC2_Wait              = 1; 
    				
    
    parameter
        wireNumPat  = 4, 
        NumRep      = 2,
        NumGsub     = 0,
        Tproj_dly   = 110,
        Tgl_res     = 200,
        Tadd        = 3,
        wireExp     = 1000,
        TLedOn      = 30000,
        Tdes2_d     = 2,
        Tdes2_w     = 4,
        Tmsken_d    = 4,
        Tmsken_w    = 11,
        Tgsub_w     = 100,
        TExpRst     = 100,
        TdrainR_d   = 10,
        TdrainF_d   = 20,
        T_MU_wait   = 1024;

    
    parameter 
    	T_DEC_SEL_0 = 2,
        T_DEC_SEL_1 = 0,
        T_DEC_EN_0  = 4,
        T_DEC_EN_1  = 0,
        T_DONE_1    = 2;

    parameter
    	TrigNo      = 1,     
        TrigOffTime = 1,            
        TrigOnTime  = 3142,
        TrigWaitTime = 100;    
    

   
    //EXP-------------------------------------- 
    Exposure_v1_T7 exposure_inst (
    	.rst(wirerst[0]),
        .CLKM(CLKMi),
    	.trigger_o(ex_trigger),
    	.re_busy(re_busy),
    	.PIXGSUBC(PIX_GSUBC),
    	.PIXDRAIN(PIX_DRAIN),
    	.PIXGLOB_RES(PIXGLOB_RES_i),
    	//.PIXGLOB_RES(PIXGLOB_RES),
    	.PIXVTG_GLOB(PIXVTG_GLOB),
    	.MASK_EN(MASK_EN),
    	.EN_STREAM(rd_enable),
    	.DES_2ND(DES2ND),
    	.PROJ_TRG(PROJ_TRG),
    	.ROWADD(ROWADD_EXP),
    	.contrastLED(contrastLED),

    	.NUM_PAT(wireNumPat),
    	.NUM_REP(NumRep),
    	.NUM_ROW(NUM_ROW),
    	.NUM_GSUB(NumGsub),
    	.Tproj_dly(Tproj_dly),
    	.Tgl_res(Tgl_res),
    	.Tadd(Tadd),
    	.Texp_ctrl(wireExp),
    	.Tdes2_d(Tdes2_d),
    	.Tdes2_w(Tdes2_w),
    	.Tmsken_d(Tmsken_d),
    	.Tmsken_w(Tmsken_w),
    	.Tgsub_w(Tgsub_w),
    	.Treset(TExpRst),
    	.TdrainR_d(TdrainR_d),
    	.TdrainF_d(TdrainF_d),
    	.T_MU_wait(T_MU_wait)
    );


    iamTriggered triggerMe(
        .clk(TX_CLKi),                      // input clk                     
        .trig_in(~PIXGLOB_RES_i),              // proj_trg generated by exposure
        .trig_out(trig_out),            // output trigger        
        .TrigNo(TrigNo),                // Number of triggers     
        .TrigOffTime(TrigOffTime),      // Off time for trigger            
        .TrigOnTime(TrigOnTime),         // On time for trigger
        .TrigWaitTime(TrigWaitTime)      // Wait time for trigger               
    );

    //wire [31:0] RO_Tcolumn_t7, RO_T1_t7, RO_T2_t7, RO_T3_t7, RO_T4_t7, RO_T5_t7, RO_T6_t7, RO_T7_t7, RO_T8_t7, RO_Treset_t7; 
    wire [8:0] ROWADD_RO_t7;
    Readout_Merge	u_Readout_Merge(
    	.rst				(wirerst[0]),
    	
    	.adc1_start_trigger (adc1_start_trigger),
    	.adc1_busy 			(adc1_busy),

    	.adc2_start_trigger (adc2_start_trigger),
    	.adc2_busy 			(adc2_busy),
    	
    	.TX_CLK				(TX_CLKi),
    	.TX_CLKx2			(TX_CLKi2),

    	.ROWADD				(ROWADD_RO_t7),
    	.SET_ROW			(SET_ROW_RO),
    	.SET_ROW_DONE 		(SET_ROW_DONE_RO | 1),

    	.PIXLEFTBUCK_SEL	(PIX_LEFTBUCK_SEL_t7),
    	.ODDCOL_EN			(ODDCOL_EN_t7),
    	.PRECH_COL			(COL_PRECH_12_t7),
    	.ADC_RST			(ADC_RST_t7),
    	.ADC_CLK			(ADC_CLK_out_t7),

    	.RST_BAR_LTCHD		(RST_BAR_LTCHD_t7),
    	.LOAD_IN			(LOAD_IN_t7),
    	.ADC_DATA_VALID		(ADC_DATA_VALID_t7),

    	.PIXREAD_SEL		(PIXREAD_SEL_t7),
    	.ADC_BIAS_EN		(ADC_BIAS_EN_t7),
    	.COLL_EN			(COLL_EN_t7),
    	.PIXRES				(PIXRES_t7),
    	
    	.ADC1_Tcolumn   	(ADC1_Tcolumn),
    	.ADC1_T1        	(ADC1_T1),
    	.ADC1_T2_1      	(ADC1_T2_1),
    	.ADC1_T2_0      	(ADC1_T2_0),
    	.ADC1_T3        	(ADC1_T3),
    	.ADC1_T4        	(ADC1_T4),
    	.ADC1_T5        	(ADC1_T5),
    	.ADC1_T6        	(ADC1_T6),   
    	.ADC1_T7        	(ADC1_T7),
    	.ADC1_T8        	(ADC1_T8),
    	.ADC1_T9        	(ADC1_T9),
    	.ADC1_TADC      	(ADC1_TADC),
    	.ADC1_NUM_ROW   	(ADC1_NUM_ROW),
    	.ADC1_Wait      	(ADC1_Wait),

    	.ADC2_Tcolumn   	(ADC2_Tcolumn),
    	.ADC2_T1        	(ADC2_T1),
    	.ADC2_T2_1      	(ADC2_T2_1),
    	.ADC2_T2_0      	(ADC2_T2_0),
    	.ADC2_T3        	(ADC2_T3),
    	.ADC2_T4        	(ADC2_T4),
    	.ADC2_T5        	(ADC2_T5),
    	.ADC2_T6        	(ADC2_T6),
    	.ADC2_T7        	(ADC2_T7),
    	.ADC2_T8        	(ADC2_T8),
    	.ADC2_T9        	(ADC2_T9),
    	.ADC2_TADC      	(ADC2_TADC),
    	.ADC2_NUM_ROW   	(ADC2_NUM_ROW),
    	.ADC2_Wait      	(ADC2_Wait)			
    );



    wire [17:1] DIGOUT;
    DIGOUT_test u_DIGOUT_test(
    	.clk			(TX_CLKi),
    	.rst			(adc2_start_trigger || adc1_start_trigger),
    	.RST_BAR_LTCHD	(RST_BAR_LTCHD_t7),
    	.ADC_DATA_VALID	(ADC_DATA_VALID),
    	.DIGOUT			(DIGOUT[17:1])
    );

    	
    ADCtoFIFO i_adc_fifo(
        .rst(wirerst[0]),
//        .adc_clk0_i(TXCLK_OUT),
        .adc_clk0_i(TX_CLKi),
        .adc_gr0_valid(ADC_DATA_VALID),
//        .adc_gr0_valid(1),
        .ch_data_i(DIGOUT[17:1]),
        .p0_rd_clk(TX_CLKi),
        .p0_rd_en(1),
        .p0_rd_data_cnt(pipe0_in_rd_count),
        .p0_full(pipe0_in_full),
        .p0_empty(pipe0_in_empty),
        .p0_valid(pipe0_in_valid),
        .p0_data_o(pipe0_in_rd_data)
    );

	assign ROWADD_RO[8:0] = adc1_busy ? ROWADD_RO_t7[8:0] : ROWADD_ADC2_MAPPED;
    wire [9:0] ROWADD_DEC;
    set_row_decoder exp_ro_row_decoder(
    	.clk(TX_CLKi),
    	.rst(wirerst[0]),

    	.ROWADD_MU(ROWADD_EXP),
    	.ROWADD_RO(ROWADD_RO[9:0]),
    	.SET_ROW_MU(DES2ND),
    	.SET_ROW_RO(SET_ROW_RO),
    
    	.SET_ROW_DONE_MU(SET_ROW_DONE_MU),
    	.SET_ROW_DONE_RO(SET_ROW_DONE_RO),
    	.DEC_SEL(DEC_SEL),     
    	.DEC_EN(DEC_EN),      
    	.ROWADD_op(ROWADD_DEC[9:0]),    
    
    	.T_DEC_SEL_0(T_DEC_SEL_0[31:0]),
    	.T_DEC_SEL_1(T_DEC_SEL_1[31:0]),
    	.T_DEC_EN_0(T_DEC_EN_0[31:0]), 
    	.T_DEC_EN_1(T_DEC_EN_1[31:0]), 
    	.T_DONE_1(T_DONE_1[31:0])    	
    );
	wire [8:0] ROWADD_ADC2_MAPPED, mem_write_addr, mem_write_data;
	row_map_table map_rows_adc2(
		.clk(TX_CLKi),
		.rowadd_in(ROWADD_RO_t7[8:0]),
		.rowadd_out(ROWADD_ADC2_MAPPED[8:0]),
		
		.mem_write_addr(mem_write_addr[8:0]), // address to write
		.mem_write_data(mem_write_data[8:0]), // what to write
		.we(0)					  // when to write
	);
  
//	assign ROWADD = (re_busy) ? ROWADD_RO : ROWADD_EXP;
    assign ROWADD = ROWADD_DEC;
    
    assign adc1_start_trigger = ex_trigger	         ;
    assign adc2_start_trigger = trig_out             ;
    
    
    assign re_busy            = adc1_busy            ;
    assign ROWADD_RO          = ROWADD_RO_t7         ;
    assign PIXREAD_EN         = PIXREAD_SEL_t7       ;
    assign PIX_LEFTBUCK_SEL   = PIX_LEFTBUCK_SEL_t7  ;
    assign PIX_RIGHTBUCK_SEL  = PIX_LEFTBUCK_SEL_t7  ;
    assign COL_PRECH_12       = COL_PRECH_12_t7      ;
    assign COLL_EN            = COLL_EN_t7           ;
    assign ODDCOL_EN          = ODDCOL_EN_t7         ;
    assign LOAD_IN            = LOAD_IN_t7           ;
    assign ADC_RST            = ADC_RST_t7           ;
    assign ADC_DATA_VALID     = ADC_DATA_VALID_t7    ;
    
    //set initial values
        integer cnt_busy = 0;
    always @(posedge clk_100) begin
    	if (rst) begin
    		//ex_trigger <= 1'b0;
    		cnt_busy <= cnt_busy + 1;
    		if (cnt_busy >= 20) begin
    		     rst <= 1'b0;
    		     cnt_busy <= 1'b0;
    		end
    	end 
    end

    //set initial values	
    initial begin
    		Select[31:0] = 32'h00000000;
    		wirerst[0] = 1;		
    #20		wirerst[0] = 0;
    
    
    end

  
endmodule
