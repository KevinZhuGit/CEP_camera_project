`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 08/18/2022 12:48:50 AM
// Design Name: 
// Module Name: iamTriggered
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module iamTriggered(
    input wire clk,                 // input clk
	input wire trig_in,             // proj_trg generated by exposure
	input wire [31:0] TrigOffTime,  // Off time for trigger
	input wire [31:0] TrigOnTime,   // On time for triggers
	input wire [31:0] TrigNo,       // Number of triggers
	input wire [31:0] TrigWaitTime, // delay time before first trigger
	output reg trig_out             // output trigger
	);
	//  Instantiation 
	/*
	iamTriggered triggerMe(
	    .clk(clk),                      // input clk                     
	    .trig_in(trig_in),              // proj_trg generated by exposure
	    .trig_out(trig_out),            // output trigger        
	    .TrigNo(TrigNo),                // Number of triggers     
	    .TrigOffTime(TrigOffTime),      // Off time for trigger
	    .TrigOnTime(TrigOnTime),         // On time for trigger                
	    .TrigWaitTime(TrigWaitTime)      // delay time before first trigger               
	);
	*/
	localparam s_idle   = 32'b1<<0;
	localparam s_wait   = 32'b1<<1; 
	localparam s_on     = 32'b1<<2;
	localparam s_off    = 32'b1<<3;
	
	integer cnt_trig    = 0;
	integer cnt_trigNo  = 0;
	integer state       = 0;
	
	reg trigReg, trigOld=0;
	
	always @ (posedge clk) begin
		case(state)
			s_idle: begin
				trigOld  <= trig_in;
				trig_out <= 0;
				state    <= trig_in && ~trigOld ? s_wait : s_idle;                        // Start only on positive edge when input trigger is asserted
				cnt_trig <= 0;                                                          // reset the counter
				cnt_trigNo <= 0;                                                        // reset the projection trigger number
			end
			s_wait: begin
				trig_out    <= 0;                                                       	// wait to assert the output trigger
				state       <= (cnt_trig == TrigWaitTime-1) ? s_on         : s_wait;         // change state after certain number of clk cycles
				cnt_trig    <= (cnt_trig == TrigWaitTime-1) ? 0            : cnt_trig + 1; // count projector Wait time
				cnt_trigNo <= 0;                                                        // reset the projection trigger number
			end
			s_on: begin
				trig_out    <= 1;                                                       // assert the output trigger
				state       <= (cnt_trig == TrigOnTime-1) ? s_off         : s_on;         // change state after certain number of clk cycles
				cnt_trig    <= (cnt_trig == TrigOnTime-1) ? 0             : cnt_trig + 1; // count projector ON time
				cnt_trigNo  <= (cnt_trig == TrigOnTime-1) ? cnt_trigNo + 1: cnt_trigNo;   // counter number of projector triggers
			end
			s_off: begin
				trig_out    <= 0;                                                                                       // de-assert the output trigger
				state       <= (cnt_trig == TrigOffTime)? ((cnt_trigNo == TrigNo) ? s_idle : s_on) : s_off;        // change state to on or idle
				cnt_trig    <= (cnt_trig == TrigOffTime) ? 0                                       : cnt_trig + 1; // count projector OFF time
			end
			default: begin
				trig_out    <= 0;
				state       <= s_idle;
				cnt_trig    <= 0;
				cnt_trigNo  <= 0;
			end
		endcase
	end

endmodule

