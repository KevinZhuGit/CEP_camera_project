`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 08/12/2020 05:33:13 PM
// Design Name: 
// Module Name: tb_proj_ctl
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module tb_proj_ctl(

    );
    

    reg clk_200,clk_25, trig_in;
    wire trig_out;
    reg [31:0] trigNo, projOnTime, projOffTime;


	reg clk_100; initial clk_100 = 1'b0; always #5   clk_100 = ~clk_100; 
	reg clk_200; initial clk_200 = 1'b0; always #2.5 clk_200 = ~clk_200; 
    reg clk_7  ; initial clk_7   = 1'b0; always #35  clk_7   = ~clk_7; 
	reg clk_25;  initial clk_25  = 1'b0; always #20   clk_25 = ~clk_25;

    wire CLKMi, TX_CLKi, TX_CLKi2;
    assign CLKMi = clk_100;
    assign TX_CLKi  = clk_100;
    assign TX_CLKi2 = clk_200;
    assign ADC_CLK  = clk_7;
	reg rst;

	wire [7:0] ROWADD;
	wire [7:0] ROWADD_EXP;
	wire [7:0] ROWADD_RO;
    
	wire ex_trigger;	
	wire re_busy;


	//RO----------------------------------------
	
	parameter
		NUM_SAMP	= 2,
		NUM_ROW		= 4,
		T_PIX		= 100,
		T1         = 5,
		T2         = 100,
		T3         = 20,
		T4         = 10,
		T5         = 14,
		T6         = 6,
		T7         = 17,
		T8         = 14,
	    TADC       = 13,
	    TOSR       = 115,
	    TReadRst   = 100,
	    Tbuck      = 1652;

    parameter
        wireNumPat  = 4,
        NumRep      = 10,
        NumGsub     = 0,
        Tproj_dly   = 38000,
        Tgl_res     = 200,
        Tadd        = 3,
//        wireExp     = 40000,
        wireExp     = 672350,
        TLedOn      = 30000,
        Tdes2_d     = 2,
        Tdes2_w     = 4,
        Tmsken_d    = 3,
        Tmsken_w    = 4,
        Tgsub_w     = 100,
        TExpRst     = 19010,
        TdrainR_d   = 10,
        TdrainF_d   = 15;
    

Readout_v1_T4	#(.NUM_ROW(10))
    u_readout_v1_T4(
	.rst(rst),
	.trigger_i(ex_trigger),
	.re_busy(re_busy),
  	.ROWADD(ROWADD_RO),
	.PIXREAD_SEL(PIXREAD_EN),
 	.PIXLEFTBUCK_SEL(PIXLEFTBUCK_SEL_i),
  	.PIXRES(PIXRES),
 	.COLLOAD_EN(),
  	.PRECH_COL(COL_PRECH),
  	//.ADC_EN_N(ADC_EN_PRE),
	.ADC_EN_N(),
  	.DATA_LOAD(DATA_LOAD),
  	.RST_ADC(RST_ADC),
 	.RST_OUTMUX(RST_OUTMUX),
  	.ADC_CLK(ADC_CLK),
	.ADC_DATA_VALID(ADC_DATA_VALID),
  	.TX_CLK(TX_CLKi),
  	.TX_CLKx2(TX_CLKi2),
	.TX_CLK_OUT(TXCLK_OUT),
//	.TX_CLK_OUT(1),
	.Tbuck(Tbuck),
	.T1(T1),
	.T2(T2),
	.T3(T3),
	.T4(T4),
	.T5(T5),
	.T6(T6),
	.T7(T7),
	.T8(T8),
	.T_ADC(TADC),
	.T_OSR(TOSR),
	.Treset(TReadRst)
    );

    
	//EXP-------------------------------------- 
    wire PIXGLOB_RES;
	Exposure_v1_T4	#(.NUM_ROW(320))
	 exposure_inst (
		.rst(rst),
        .CLKM(CLKMi),
		.trigger_o(ex_trigger),
		.re_busy(re_busy),
		.PIXGSUBC(PIXGSUBC),
		.PIXDRAIN(PIXDRAIN),
//		.PIXGLOB_RES(PIXGLOB_RES_i),
		.PIXGLOB_RES(PIXGLOB_RES),
		.PIXVTG_GLOB(PIXVTG_GLOB),
		.MASK_EN(MASK_EN),
		.EN_STREAM(rd_enable),
		.DES_2ND(DES),
		.PROJ_TRG(PROJ_TRG),
		.ROWADD(ROWADD_EXP),
		.contrastLED(contrastLED),

		.NUM_PAT(wireNumPat),
		.NUM_REP(NumRep),
		.NUM_GSUB(NumGsub),
		.Tproj_dly(Tproj_dly),
		.Tgl_res(Tgl_res),
		.Tadd(Tadd),
		.Texp_ctrl(wireExp),
		.Tdes2_d(Tdes2_d),
		.Tdes2_w(Tdes2_w),
		.Tmsken_d(Tmsken_d),
		.Tmsken_w(Tmsken_w),
		.Tgsub_w(Tgsub_w),
		.Treset(TExpRst),
		.TdrainR_d(TdrainR_d),
		.TdrainF_d(TdrainF_d),
	    .TLedOn(TLedOn)
	);

	assign ROWADD = (re_busy) ? ROWADD_RO : ROWADD_EXP;

	
	//set initial values
	    integer cnt_busy = 0;
    always @(posedge clk_100) begin
		if (rst) begin
			//ex_trigger <= 1'b0;
			cnt_busy <= cnt_busy + 1;
			if (cnt_busy >= 20) begin
			     rst <= 1'b0;
			     cnt_busy <= 1'b0;
			end
		end 
    end
    //set initial values
    
	initial begin
	       rst = 1'b1;
    #20	   rst = 0;
    
	end

    
    proj_ctl DUT(
        .clk(CLKMi),                  // input clk                     
        .trig_in(PROJ_TRG),              // proj_trg generated by exposure
        .trig_out(trig_out),            // Off time for projector        
        .trigNo(trigNo),                // On time for projector         
        .projOffTime(projOffTime),      // Number of triggers            
        .projOnTime(projOnTime)         // output trigger                
    );
    
    initial begin
        clk_200     = 0;
        clk_25      = 0;
        trig_in     = 0;
        trigNo      = 24;
        projOffTime = 70*1000/5;
        projOnTime  = 70*1000/5; 
    
        #200 trig_in = 1;
        #20 trig_in = 0;
    
        #4980 trig_in = 1;
        #20 trig_in = 0;
    end
	
    
endmodule
