`timescale 1ns / 1ps

module ADC_FIFO_ctrl();

    

endmodule // ADC_FIFO_ctrl